`timescale 1ns / 1ps


module REG_PIPE_4(
    input clk,
    input rst,
    input WB_EN,
    input MEM_R_EN,
    input [31:0] ALU_Res,
    input [31:0] MEM_Result,
    input [3:0]  Dest,

    output reg WB_EN_out,
    output reg MEM_R_EN_out,
    output reg [31:0] ALU_Res_out,
    output reg [31:0] MEM_Result_out,
    output reg [3:0]  Dest_out,
);
    
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            WB_EN_out <= 1'b0;
            MEM_R_EN_out <= 1'b0;
            ALU_Res_out <= 32'b0;
            MEM_Result_out <= 32'b0;
            Dest_out <= 4'b0;
        end else begin
            WB_EN_out <= WB_EN;
            MEM_R_EN_out <= MEM_R_EN;
            ALU_Res_out <= ALU_Res;
            MEM_Result_out <= MEM_Result;
            Dest_out <= Dest;
        end
    end
    
endmodule