`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/20/2025 04:38:18 PM
// Design Name: 
// Module Name: EX_stage
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module EXE_STAGE(
    input clk,
    input rst,
    input [31:0] pc,
    input [31:0] instruction_memory,
    output wire flush,
    output reg [31:0] output_pc,
    output reg [31:0] output_instruction_memory
);
    
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            output_pc <= 32'b0;
            output_instruction_memory <= 32'b0;
        end else begin
            // Normal operation
            output_pc <= pc;
            output_instruction_memory <= instruction_memory;
        end
    end
    assign flush = 0;
    
endmodule